library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- entity combinational including 3 inputs and 1 output -- 
entity combinational is
	PORT( a, b, c : in STD_LOGIC;
			f : out STD_LOGIC
			);
end combinational;


-- behaviour of the combinational circuit -- 
architecture Behavioural of combinational is
begin
	f <= (((NOT a) AND b) OR ((NOT A) AND c) OR ((NOT b) OR c) OR (a OR (NOT b))); -- assign equation to f -- 
end Behavioural;

