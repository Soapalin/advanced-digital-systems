library IEEE;
use IEEE.STD-LOGIC-1164.ALL;

entity stringcheck is 
	PORT(
		input: IN STD_LOGIC;
		output: OUT STD_LOGIC
		);
end stringcheck;



architecture behaviour of stringcheck is 
BEGIN



END behaviour;